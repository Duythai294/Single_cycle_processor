`timescale 1ns / 1ps

module Mux_tb;

    // Inputs
    reg [31:0] a, b;
    reg s;

    // Output
    wire [31:0] c;

    Mux uut (
        .a(a),
        .b(b),
        .s(s),
        .c(c)
    );

    initial begin
        $display("----- Mux Testbench -----");
        
        // Test 1: s = 0 => output = a
        a = 32'hAAAAAAAA;
        b = 32'h55555555;
        s = 0;
        #10;
        $display("s=%b | a=0x%h | b=0x%h | c=0x%h (Expect a)", s, a, b, c);

        // Test 2: s = 1 => output = b
        s = 1;
        #10;
        $display("s=%b | a=0x%h | b=0x%h | c=0x%h (Expect b)", s, a, b, c);

        // Test 3: a = 0, b = 0xFFFFFFFF, s = 0 => expect a
        a = 32'h00000000;
        b = 32'hFFFFFFFF;
        s = 0;
        #10;
        $display("s=%b | a=0x%h | b=0x%h | c=0x%h (Expect a)", s, a, b, c);

        // Test 4: s = 1 => expect b
        s = 1;
        #10;
        $display("s=%b | a=0x%h | b=0x%h | c=0x%h (Expect b)", s, a, b, c);

        $finish;
    end

endmodule

